-- Bus functional model
-- $URL: $
