-- Top-level
-- $URL $
