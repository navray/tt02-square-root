-- Top-level
-- $URL: $
